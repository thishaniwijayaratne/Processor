module IRAM(input clk,
				input [6:0] PC,
				output reg [19:0] instr_out);
				
	reg [19:0] ram [44:0];	//Needs to change
	
//	parameter = 

	
	initial begin
		ram [0]  = 0011 000000000000 0001; //write 0000 Ax;
		ram [1]  = 0011 010000000000 0010; //write 1024 Ay
		ram [2]  = 0011 100000000000 0011; //write 2048 Az
		
		ram [3]  = 0100 110000000000 0100; //LOADI 3072 Rx
		ram [4]  = 0100 110000000001 0101; //LOADI 3073 Cx
		ram [5]  = 0100 110000000010 0110; //LOADI 3074 Cy
		
		ram [6]  = 0101 0101 0110 00000000 ; //MUL Cx Cy
		
		ram [7]  = 0111 1110 000000000000; //MV Sy
		
		ram [8]  = 0010 1000 000000000000; //RST TR2
		ram [9]  = 0010 1011 000000000000; //RST I
		ram [10] = 0010 1100 000000000000; //RST J
		ram [11] = 0010 1101 000000000000; //RST K
		
		ram [12] = 0110 1001 0001 00000000; //LOAD Vx Ax
		ram [13] = 0110 1010 0010 00000000; //LOAD Vy Ay
		ram [14] = 0101 1001 1010 00000000; //MUL Vx Vy
		ram [15] = 0111 0111 000000000000; //MV TR1
		ram [16] = 1000 0111 1000 00000000; //ADD TR1 TR2
		ram [17] = 0111 1000 000000000000; //MV TR2
		
		ram [18] = 1001 1101 000000000000; //INC K
		ram [19] = 1010 0101 1101 00000000; //SUB Cx K
		ram [20] = 1011 100001 0000000000; //JMPZ 33
		
		//Jumped..............
		
		ram [21] = 0010 1101 000000000000; //RST K		
		ram [22] = 1101 1000 0011 00000000 ; //STORE TR2 Az
		ram [23] = 1001 0011 000000000000; //INC Az
		
		ram [24] = 0010 1000 000000000000; //RST TR2
		ram [25] = 1001 1100 000000000000; //INC J
		ram [26] = 1010 0110 1100 00000000; //SUB Cy J
		ram [27] = 1011 100100 0000000000; //JUMPZ 36
		
		ram [28] = 0010 1100 000000000000; //RST J
		ram [29] = 1001 1011 000000000000; //INC I	
		ram [30] = 1010 0100 1010 00000000; //SUB Rx I
		ram [31] = 1011 101001 0000000000; //JUMPZ 41
		ram [32] = 1110 000000000000 0000; //END ?????????????????????????????????????????????????????
		

		ram [33] = 1001 0001 000000000000; //INC Ax
		ram [34] = 1001 0010 000000000000; //INC Ay
		ram [35] = 1100 001100 0000000000; //JMP 12
		
		ram [36] = 1001 0010 000000000000; //INC Ay
		ram [37] = 1001 0001 000000000000; //INC Ax
		ram [38] = 1010 0001 0101 00000000; //SUB Ax Cx
		ram [39] = 0111 0001 000000000000; //MV Ax
		ram [40] = 1100 001100 0000000000; //JMP 12
		
		
		ram [41] = 1001 0001 000000000000; //INC Ax
		ram [42] = 1001 0010 000000000000; //INC Ay
		ram [43] = 1010 0010 1110 00000000; //SUB Ay Sy
		ram [44] = 0111 0010 000000000000; //MV Ay
		ram [45] = 1100 001100 0000000000; //JMP 12
	
	end
	
	
	always @(posedge clk)begin
		instr_out = ram[PC];		
		
	end
	

endmodule 