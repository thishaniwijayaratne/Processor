module Input_data();

endmodule