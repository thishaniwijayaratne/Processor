module DRAM();

endmodule