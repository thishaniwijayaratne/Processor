module Store_data();

endmodule