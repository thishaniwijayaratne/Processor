module IRAM(input clk,
				input [5:0] PC,
				output reg [19:0] instr_out);
				
	reg [19:0] ram [44:0];	//Needs to change
	
	initial begin
		ram [0]  = 00110001000000000000; //write Ax 0000;
		ram [1]  = 00110010010000000000; //write Ay 1024 
		ram [2]  = 00110011100000000000; //write Az 2048 
		
		ram [3]  = 01000100110000000000; //LOADI 3072 Rx
		ram [4]  = 01000101110000000001; //LOADI 3073 Cx
		ram [5]  = 01000110110000000010; //LOADI 3074 Cy
		
		ram [6]  = 01010101011000000000; //MUL Cx Cy
		
		ram [7]  = 01111110000000000000; //MV Sy
		
		ram [8]  = 00101000000000000000; //RST TR2
		ram [9]  = 00101011000000000000; //RST I
		ram [10] = 00101100000000000000; //RST J
		ram [11] = 00101101000000000000; //RST K
		
		ram [12] = 01101001000100000000; //LOAD Vx Ax
		ram [13] = 01101010001000000000; //LOAD Vy Ay
		ram [14] = 01011001101000000000; //MUL Vx Vy
		ram [15] = 01110111000000000000; //MV TR1
		ram [16] = 10000111100000000000; //ADD TR1 TR2
		ram [17] = 01111000000000000000; //MV TR2
		
		ram [18] = 10011101000000000000; //INC K
		ram [19] = 10100101110100000000; //SUB Cx K
		ram [20] = 10111000010000000000; //JMPZ 33
		
		//Jumped..............
		
		ram [21] = 00101101000000000000; //RST K		
		ram [22] = 11011000001100000000; //STORE TR2 Az
		ram [23] = 10010011000000000000; //INC Az
		
		ram [24] = 00101000000000000000; //RST TR2
		ram [25] = 10011100000000000000; //INC J
		ram [26] = 10100110110000000000; //SUB Cy J
		ram [27] = 10111001000000000000; //JUMPZ 36
		
		ram [28] = 00101100000000000000; //RST J
		ram [29] = 10011011000000000000; //INC I	
		ram [30] = 10100100101000000000; //SUB Rx I
		ram [31] = 10111010010000000000; //JUMPZ 41
		ram [32] = 11100000000000000000; //END ?????????????????????????????????????????????????????
		

		ram [33] = 10010001000000000000; //INC Ax
		ram [34] = 10010010000000000000; //INC Ay
		ram [35] = 11000011000000000000; //JMP 12
		
		ram [36] = 10010010000000000000; //INC Ay
		ram [37] = 10010001000000000000; //INC Ax
		ram [38] = 10100001010100000000; //SUB Ax Cx
		ram [39] = 01110001000000000000; //MV Ax
		ram [40] = 11000011000000000000; //JMP 12
		
		
		ram [41] = 10010001000000000000; //INC Ax
		ram [42] = 10010010000000000000; //INC Ay
		ram [43] = 10100010111000000000; //SUB Ay Sy
		ram [44] = 01110010000000000000; //MV Ay
		ram [45] = 11000011000000000000; //JMP 12
	
	end
	
	
	always @(posedge clk)begin
		instr_out = ram[PC];		
		
	end
	

endmodule 